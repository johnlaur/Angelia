// megafunction wizard: %LPM_MULT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_mult 

// ============================================================
// File Name: mult_24Sx24S.v
// Megafunction Name(s):
// 			lpm_mult
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 11.1 Build 259 01/25/2012 SP 2 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module mult_24Sx24S (
	aclr,
	clock,
	dataa,
	datab,
	result);

	input	  aclr;
	input	  clock;
	input	[23:0]  dataa;
	input	[23:0]  datab;
	output	[47:0]  result;

	wire [47:0] sub_wire0;
	wire [47:0] result = sub_wire0[47:0];

	lpm_mult	lpm_mult_component (
				.aclr (aclr),
				.clock (clock),
				.datab (datab),
				.dataa (dataa),
				.result (sub_wire0),
				.clken (1'b1),
				.sum (1'b0));
	defparam
		lpm_mult_component.lpm_hint = "MAXIMIZE_SPEED=9",
		lpm_mult_component.lpm_pipeline = 3,
		lpm_mult_component.lpm_representation = "SIGNED",
		lpm_mult_component.lpm_type = "LPM_MULT",
		lpm_mult_component.lpm_widtha = 24,
		lpm_mult_component.lpm_widthb = 24,
		lpm_mult_component.lpm_widthp = 48;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: AutoSizeResult NUMERIC "1"
// Retrieval info: PRIVATE: B_isConstant NUMERIC "0"
// Retrieval info: PRIVATE: ConstantB NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "3"
// Retrieval info: PRIVATE: Latency NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: SignedMult NUMERIC "1"
// Retrieval info: PRIVATE: USE_MULT NUMERIC "1"
// Retrieval info: PRIVATE: ValidConstant NUMERIC "0"
// Retrieval info: PRIVATE: WidthA NUMERIC "24"
// Retrieval info: PRIVATE: WidthB NUMERIC "24"
// Retrieval info: PRIVATE: WidthP NUMERIC "48"
// Retrieval info: PRIVATE: aclr NUMERIC "1"
// Retrieval info: PRIVATE: clken NUMERIC "0"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: PRIVATE: optimize NUMERIC "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_HINT STRING "MAXIMIZE_SPEED=9"
// Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "3"
// Retrieval info: CONSTANT: LPM_REPRESENTATION STRING "SIGNED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MULT"
// Retrieval info: CONSTANT: LPM_WIDTHA NUMERIC "24"
// Retrieval info: CONSTANT: LPM_WIDTHB NUMERIC "24"
// Retrieval info: CONSTANT: LPM_WIDTHP NUMERIC "48"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL "aclr"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: dataa 0 0 24 0 INPUT NODEFVAL "dataa[23..0]"
// Retrieval info: USED_PORT: datab 0 0 24 0 INPUT NODEFVAL "datab[23..0]"
// Retrieval info: USED_PORT: result 0 0 48 0 OUTPUT NODEFVAL "result[47..0]"
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @dataa 0 0 24 0 dataa 0 0 24 0
// Retrieval info: CONNECT: @datab 0 0 24 0 datab 0 0 24 0
// Retrieval info: CONNECT: result 0 0 48 0 @result 0 0 48 0
// Retrieval info: GEN_FILE: TYPE_NORMAL mult_24Sx24S.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult_24Sx24S.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult_24Sx24S.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult_24Sx24S.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult_24Sx24S_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult_24Sx24S_bb.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult_24Sx24S_waveforms.html FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mult_24Sx24S_wave*.jpg FALSE
// Retrieval info: LIB_FILE: lpm
